-- Ryan Raghani – 301623888; Danny Woo – 301613129; Mitchell Kieper – 301590274;


-- second part of the package file to declare direction_t
library ieee;
use ieee.std_logic_1164.all;

package body elevator_types is
end package body elevator_types;
