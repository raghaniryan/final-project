-- Ryan Raghani – 301623888; Danny Woo – 301613129; Mitchell Kieper – 301590274;


-- no longer used in the project
